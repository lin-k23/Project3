.title testbench for muxiplexer
.include "..\simlib.sp"

* ########################Multiplexer model######################## *
.subckt muxiplexer A B S Z VDD VSS
.ends muxiplexer