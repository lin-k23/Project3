.title testbench for Full Adder
.include "..\simlib.sp"

.subckt FA A B C Z VDD VSS
* ########################Full Adder model######################## *

.ends FA